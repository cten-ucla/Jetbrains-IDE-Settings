Title
*==============================================================================


.end